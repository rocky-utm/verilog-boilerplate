module NAME();
// definition
endmodule

module NAME_tb();
//definitions

NAME NAME_inst(
//map
);

initial begin
//process
end
endmodule
